`include "uvm_macros.svh"
import uvm_pkg::*;

class dut_agent extends uvm_agent;

  `uvm_component_utils(dut_agent)

  uvm_sequencer #(dut_txn) seqr;
  dut_driver  drv;
  dut_monitor mon;

  // ✅ REQUIRED constructor
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    seqr = uvm_sequencer #(dut_txn)::type_id::create("seqr", this);
    drv  = dut_driver ::type_id::create("drv",  this);
    mon  = dut_monitor::type_id::create("mon",  this);
  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    drv.seq_item_port.connect(seqr.seq_item_export);
  endfunction

endclass